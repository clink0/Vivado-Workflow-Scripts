module SSDispFLC(clk, seg, dp, an);
input clk;
output dp;
output reg [6:0] seg;
output reg [3:0] an;

reg [1:0] state = 2'b00;
assign dp = 1'b1;
parameter cntmax = 10'd1023;
reg [9:0] cnt;

always @(posedge clk)
begin
  if(cnt == cntmax)
  begin
    if (state == 2'b00)
       begin
         cnt <= 0;
	 an <= 4'b1110;
	 seg <= 7'b1000110;
	 state <= state + 1;
       end

    else if (state == 2'b01)
       begin
         cnt <= 0;
	 an <= 4'b1101;
	 seg <= 7'b1000111;
	 state <= state + 1;
       end

    else if (state == 2'b10)
       begin
         cnt <= 0;
	 an <= 4'b1011;
	 seg <= 7'b0001110;
	 state <= 2'b00;
       end
  end
  else cnt <= cnt + 1;
end
endmodule
