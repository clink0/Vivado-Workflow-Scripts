module SSDisp(clk, an, seg, dp, sw);
input clk;
input [3:0] sw;
output [3:0] an;
output reg [6:0] seg;
output dp;

assign dp = 1'b1;
assign an[3:0] = 4'b1110;

always @ (posedge clk)
begin
  case(sw)
                    
  4'b0000 : seg <= 7'b1000000;
  4'b0001 : seg <= 7'b1111001;
  4'b0010 : seg <= 7'b0100100;
  4'b0011 : seg <= 7'b0110000;
  4'b0100 : seg <= 7'b0011001;
  4'b0101 : seg <= 7'b0010010;
  4'b0110 : seg <= 7'b0000010;
  4'b0111 : seg <= 7'b1111000;
  4'b1000 : seg <= 7'b0000000;
  4'b1001 : seg <= 7'b0010000;
  
  endcase

end
endmodule
